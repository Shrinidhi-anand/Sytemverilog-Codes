// Code your design here

class packet;
  rand bit [2:0]addr1;
  randc bit [2:0]addr2;
endclass