// Code your design here

