// Code your design here

class packet;
  rand bit [2:0]addr;
  randc bit [2:0]data;
endclass