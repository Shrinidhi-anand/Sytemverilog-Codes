// Code your design here


  class A;
    integer m;
  endclass